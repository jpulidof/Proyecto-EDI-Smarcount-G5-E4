// output_driver.v
// Módulo de salida SOLO con display 7 segmentos (Cyclone IV)

module output_driver (
    input wire [1:0] color_code,
    output reg [6:0] seg  // Display de 7 segmentos (activo en 0)
);

    always @(*) begin
        // Mostrar una letra en el display según el color detectado
        case (color_code)
            2'b00: seg = 7'b1000110; // 'r' (forma simplificada)
            2'b01: seg = 7'b0001000; // 'G'
            2'b10: seg = 7'b0010010; // 'b'
            default: seg = 7'b1111110; // '-' para desconocido
        endcase
    end

endmodule
